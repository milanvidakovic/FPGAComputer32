module ROM#(parameter N = 5'd16)(
    input [31:0] addr,
	 input rd,
    output reg [15:0] data
    );

always @(*)
  case (addr)

9'h000: data = 16'h0001;
9'h001: data = 16'h0000;
9'h002: data = 16'h0100;
9'h003: data = 16'h0000;
9'h004: data = 16'h0000;
9'h005: data = 16'h0000;
9'h006: data = 16'h0000;
9'h007: data = 16'h0000;
9'h008: data = 16'h0000;
9'h009: data = 16'h0000;
9'h00A: data = 16'h0000;
9'h00B: data = 16'h0000;
9'h00C: data = 16'h0000;
9'h00D: data = 16'h0000;
9'h00E: data = 16'h0000;
9'h00F: data = 16'h0000;
9'h010: data = 16'h0000;
9'h011: data = 16'h0000;
9'h012: data = 16'h0000;
9'h013: data = 16'h0000;
9'h014: data = 16'h0000;
9'h015: data = 16'h0000;
9'h016: data = 16'h0000;
9'h017: data = 16'h0000;
9'h018: data = 16'h0000;
9'h019: data = 16'h0000;
9'h01A: data = 16'h0000;
9'h01B: data = 16'h0000;
9'h01C: data = 16'h0000;
9'h01D: data = 16'h0000;
9'h01E: data = 16'h0000;
9'h01F: data = 16'h0000;
9'h020: data = 16'h0000;
9'h021: data = 16'h0000;
9'h022: data = 16'h0000;
9'h023: data = 16'h0000;
9'h024: data = 16'h0000;
9'h025: data = 16'h0000;
9'h026: data = 16'h0000;
9'h027: data = 16'h0000;
9'h028: data = 16'h0000;
9'h029: data = 16'h0000;
9'h02A: data = 16'h0000;
9'h02B: data = 16'h0000;
9'h02C: data = 16'h0000;
9'h02D: data = 16'h0000;
9'h02E: data = 16'h0000;
9'h02F: data = 16'h0000;
9'h030: data = 16'h0000;
9'h031: data = 16'h0000;
9'h032: data = 16'h0000;
9'h033: data = 16'h0000;
9'h034: data = 16'h0000;
9'h035: data = 16'h0000;
9'h036: data = 16'h0000;
9'h037: data = 16'h0000;
9'h038: data = 16'h0000;
9'h039: data = 16'h0000;
9'h03A: data = 16'h0000;
9'h03B: data = 16'h0000;
9'h03C: data = 16'h0000;
9'h03D: data = 16'h0000;
9'h03E: data = 16'h0000;
9'h03F: data = 16'h0000;
9'h040: data = 16'h0000;
9'h041: data = 16'h0000;
9'h042: data = 16'h0000;
9'h043: data = 16'h0000;
9'h044: data = 16'h0000;
9'h045: data = 16'h0000;
9'h046: data = 16'h0000;
9'h047: data = 16'h0000;
9'h048: data = 16'h0000;
9'h049: data = 16'h0000;
9'h04A: data = 16'h0000;
9'h04B: data = 16'h0000;
9'h04C: data = 16'h0000;
9'h04D: data = 16'h0000;
9'h04E: data = 16'h0000;
9'h04F: data = 16'h0000;
9'h050: data = 16'h0000;
9'h051: data = 16'h0000;
9'h052: data = 16'h0000;
9'h053: data = 16'h0000;
9'h054: data = 16'h0000;
9'h055: data = 16'h0000;
9'h056: data = 16'h0000;
9'h057: data = 16'h0000;
9'h058: data = 16'h0000;
9'h059: data = 16'h0000;
9'h05A: data = 16'h0000;
9'h05B: data = 16'h0000;
9'h05C: data = 16'h0000;
9'h05D: data = 16'h0000;
9'h05E: data = 16'h0000;
9'h05F: data = 16'h0000;
9'h060: data = 16'h0000;
9'h061: data = 16'h0000;
9'h062: data = 16'h0000;
9'h063: data = 16'h0000;
9'h064: data = 16'h0000;
9'h065: data = 16'h0000;
9'h066: data = 16'h0000;
9'h067: data = 16'h0000;
9'h068: data = 16'h0000;
9'h069: data = 16'h0000;
9'h06A: data = 16'h0000;
9'h06B: data = 16'h0000;
9'h06C: data = 16'h0000;
9'h06D: data = 16'h0000;
9'h06E: data = 16'h0000;
9'h06F: data = 16'h0000;
9'h070: data = 16'h0000;
9'h071: data = 16'h0000;
9'h072: data = 16'h0000;
9'h073: data = 16'h0000;
9'h074: data = 16'h0000;
9'h075: data = 16'h0000;
9'h076: data = 16'h0000;
9'h077: data = 16'h0000;
9'h078: data = 16'h0000;
9'h079: data = 16'h0000;
9'h07A: data = 16'h0000;
9'h07B: data = 16'h0000;
9'h07C: data = 16'h0000;
9'h07D: data = 16'h0000;
9'h07E: data = 16'h0000;
9'h07F: data = 16'h0000;
9'h080: data = 16'h0FB0;
9'h081: data = 16'h0000;
9'h082: data = 16'h3000;
9'h083: data = 16'h0020;
9'h084: data = 16'h0001;
9'h085: data = 16'h0120;
9'h086: data = 16'h0010;
9'h087: data = 16'h0183;
9'h088: data = 16'h00B0;
9'h089: data = 16'h0000;
9'h08A: data = 16'h0238;
9'h08B: data = 16'h01B0;
9'h08C: data = 16'h0000;
9'h08D: data = 16'h0012;
9'h08E: data = 16'h018C;
9'h08F: data = 16'h00B0;
9'h090: data = 16'h0000;
9'h091: data = 16'h0000;
9'h092: data = 16'h009C;
9'h093: data = 16'h0000;
9'h094: data = 16'h038A;
9'h095: data = 16'h009C;
9'h096: data = 16'h0000;
9'h097: data = 16'h038E;
9'h098: data = 16'h009C;
9'h099: data = 16'h0000;
9'h09A: data = 16'h039E;
9'h09B: data = 16'h009C;
9'h09C: data = 16'h0000;
9'h09D: data = 16'h0392;
9'h09E: data = 16'h009C;
9'h09F: data = 16'h0000;
9'h0A0: data = 16'h03A2;
9'h0A1: data = 16'h00B0;
9'h0A2: data = 16'h0000;
9'h0A3: data = 16'hB000;
9'h0A4: data = 16'h009C;
9'h0A5: data = 16'h0000;
9'h0A6: data = 16'h0396;
9'h0A7: data = 16'h0002;
9'h0A8: data = 16'h0000;
9'h0A9: data = 16'h0214;
9'h0AA: data = 16'h0002;
9'h0AB: data = 16'h0000;
9'h0AC: data = 16'h01DE;
9'h0AD: data = 16'h00B0;
9'h0AE: data = 16'h0000;
9'h0AF: data = 16'h004D;
9'h0B0: data = 16'h0002;
9'h0B1: data = 16'h0000;
9'h0B2: data = 16'h01BC;
9'h0B3: data = 16'h00B0;
9'h0B4: data = 16'h0000;
9'h0B5: data = 16'h000D;
9'h0B6: data = 16'h0002;
9'h0B7: data = 16'h0000;
9'h0B8: data = 16'h01BC;
9'h0B9: data = 16'h00B0;
9'h0BA: data = 16'h0000;
9'h0BB: data = 16'h000A;
9'h0BC: data = 16'h0002;
9'h0BD: data = 16'h0000;
9'h0BE: data = 16'h01BC;
9'h0BF: data = 16'h00B0;
9'h0C0: data = 16'h0000;
9'h0C1: data = 16'h0003;
9'h0C2: data = 16'h0002;
9'h0C3: data = 16'h0000;
9'h0C4: data = 16'h01BC;
9'h0C5: data = 16'h00B0;
9'h0C6: data = 16'h0000;
9'h0C7: data = 16'h0003;
9'h0C8: data = 16'h0002;
9'h0C9: data = 16'h0000;
9'h0CA: data = 16'h01BC;
9'h0CB: data = 16'h00B0;
9'h0CC: data = 16'h0000;
9'h0CD: data = 16'h0003;
9'h0CE: data = 16'h0002;
9'h0CF: data = 16'h0000;
9'h0D0: data = 16'h01BC;
9'h0D1: data = 16'h001C;
9'h0D2: data = 16'h0000;
9'h0D3: data = 16'h039E;
9'h0D4: data = 16'h009D;
9'h0D5: data = 16'h0000;
9'h0D6: data = 16'h0001;
9'h0D7: data = 16'h0011;
9'h0D8: data = 16'h0000;
9'h0D9: data = 16'hB000;
9'h0DA: data = 16'h0000;
9'h0DB: data = 16'h0001;
9'h0DC: data = 16'h0000;
9'h0DD: data = 16'h01A2;
9'h0DE: data = 16'h0150;
9'h0DF: data = 16'h0130;
9'h0E0: data = 16'h0041;
9'h0E1: data = 16'h019D;
9'h0E2: data = 16'h0000;
9'h0E3: data = 16'h0000;
9'h0E4: data = 16'h0011;
9'h0E5: data = 16'h0000;
9'h0E6: data = 16'h01D6;
9'h0E7: data = 16'h0000;
9'h0E8: data = 16'h0001;
9'h0E9: data = 16'h0000;
9'h0EA: data = 16'h01BE;
9'h0EB: data = 16'h0040;
9'h0EC: data = 16'h0042;
9'h0ED: data = 16'h0170;
9'h0EE: data = 16'h0080;
9'h0EF: data = 16'h02B0;
9'h0F0: data = 16'h0000;
9'h0F1: data = 16'h0400;
9'h0F2: data = 16'h01B0;
9'h0F3: data = 16'h0000;
9'h0F4: data = 16'h0208;
9'h0F5: data = 16'h1033;
9'h0F6: data = 16'h009E;
9'h0F7: data = 16'h0000;
9'h0F8: data = 16'h0011;
9'h0F9: data = 16'h0000;
9'h0FA: data = 16'h0206;
9'h0FB: data = 16'h0283;
9'h0FC: data = 16'h0109;
9'h0FD: data = 16'h020D;
9'h0FE: data = 16'h0000;
9'h0FF: data = 16'h0002;
9'h100: data = 16'h0001;
9'h101: data = 16'h0000;
9'h102: data = 16'h01EA;
9'h103: data = 16'h0080;
9'h104: data = 16'h5741;
9'h105: data = 16'h4954;
9'h106: data = 16'h494E;
9'h107: data = 16'h472E;
9'h108: data = 16'h2E2E;
9'h109: data = 16'h0000;
9'h10A: data = 16'h00B0;
9'h10B: data = 16'h0000;
9'h10C: data = 16'h0000;
9'h10D: data = 16'h01B0;
9'h10E: data = 16'h0000;
9'h10F: data = 16'h0400;
9'h110: data = 16'h02B0;
9'h111: data = 16'h0000;
9'h112: data = 16'h00F0;
9'h113: data = 16'h0183;
9'h114: data = 16'h010D;
9'h115: data = 16'h0000;
9'h116: data = 16'h0002;
9'h117: data = 16'h0289;
9'h118: data = 16'h0071;
9'h119: data = 16'h0000;
9'h11A: data = 16'h0226;
9'h11B: data = 16'h0080;
9'h11C: data = 16'h0050;
9'h11D: data = 16'h0150;
9'h11E: data = 16'h0250;
9'h11F: data = 16'h0350;
9'h120: data = 16'h001C;
9'h121: data = 16'h0000;
9'h122: data = 16'h038A;
9'h123: data = 16'h009D;
9'h124: data = 16'h0000;
9'h125: data = 16'h0000;
9'h126: data = 16'h0011;
9'h127: data = 16'h0000;
9'h128: data = 16'h02F0;
9'h129: data = 16'h009D;
9'h12A: data = 16'h0000;
9'h12B: data = 16'h0001;
9'h12C: data = 16'h0011;
9'h12D: data = 16'h0000;
9'h12E: data = 16'h030E;
9'h12F: data = 16'h009D;
9'h130: data = 16'h0000;
9'h131: data = 16'h0002;
9'h132: data = 16'h0011;
9'h133: data = 16'h0000;
9'h134: data = 16'h033A;
9'h135: data = 16'h009D;
9'h136: data = 16'h0000;
9'h137: data = 16'h0003;
9'h138: data = 16'h0011;
9'h139: data = 16'h0000;
9'h13A: data = 16'h034E;
9'h13B: data = 16'h0130;
9'h13C: data = 16'h0040;
9'h13D: data = 16'h001C;
9'h13E: data = 16'h0000;
9'h13F: data = 16'h03A2;
9'h140: data = 16'h1004;
9'h141: data = 16'h009C;
9'h142: data = 16'h0000;
9'h143: data = 16'h03A2;
9'h144: data = 16'h021C;
9'h145: data = 16'h0000;
9'h146: data = 16'h0396;
9'h147: data = 16'h12B3;
9'h148: data = 16'h0209;
9'h149: data = 16'h209C;
9'h14A: data = 16'h0000;
9'h14B: data = 16'h0396;
9'h14C: data = 16'h021C;
9'h14D: data = 16'h0000;
9'h14E: data = 16'h0392;
9'h14F: data = 16'h0209;
9'h150: data = 16'h209C;
9'h151: data = 16'h0000;
9'h152: data = 16'h0392;
9'h153: data = 16'h031C;
9'h154: data = 16'h0000;
9'h155: data = 16'h038E;
9'h156: data = 16'h320A;
9'h157: data = 16'h0011;
9'h158: data = 16'h0000;
9'h159: data = 16'h02BA;
9'h15A: data = 16'h0001;
9'h15B: data = 16'h0000;
9'h15C: data = 16'h0380;
9'h15D: data = 16'h001C;
9'h15E: data = 16'h0000;
9'h15F: data = 16'h03A2;
9'h160: data = 16'h002D;
9'h161: data = 16'h0000;
9'h162: data = 16'h00FF;
9'h163: data = 16'h0002;
9'h164: data = 16'h0000;
9'h165: data = 16'h01BC;
9'h166: data = 16'h001C;
9'h167: data = 16'h0000;
9'h168: data = 16'h03A2;
9'h169: data = 16'h006D;
9'h16A: data = 16'h0000;
9'h16B: data = 16'h0008;
9'h16C: data = 16'h0002;
9'h16D: data = 16'h0000;
9'h16E: data = 16'h01BC;
9'h16F: data = 16'h00B0;
9'h170: data = 16'h0000;
9'h171: data = 16'h0001;
9'h172: data = 16'h009C;
9'h173: data = 16'h0000;
9'h174: data = 16'h039E;
9'h175: data = 16'h0001;
9'h176: data = 16'h0000;
9'h177: data = 16'h0380;
9'h178: data = 16'h0130;
9'h179: data = 16'h0040;
9'h17A: data = 16'h109C;
9'h17B: data = 16'h0000;
9'h17C: data = 16'h038E;
9'h17D: data = 16'h011C;
9'h17E: data = 16'h0000;
9'h17F: data = 16'h038A;
9'h180: data = 16'h0109;
9'h181: data = 16'h109C;
9'h182: data = 16'h0000;
9'h183: data = 16'h038A;
9'h184: data = 16'h0001;
9'h185: data = 16'h0000;
9'h186: data = 16'h0380;
9'h187: data = 16'h0130;
9'h188: data = 16'h0040;
9'h189: data = 16'h021C;
9'h18A: data = 16'h0000;
9'h18B: data = 16'h038E;
9'h18C: data = 16'h015D;
9'h18D: data = 16'h0000;
9'h18E: data = 16'h0008;
9'h18F: data = 16'h2185;
9'h190: data = 16'h109C;
9'h191: data = 16'h0000;
9'h192: data = 16'h038E;
9'h193: data = 16'h011C;
9'h194: data = 16'h0000;
9'h195: data = 16'h038A;
9'h196: data = 16'h0109;
9'h197: data = 16'h109C;
9'h198: data = 16'h0000;
9'h199: data = 16'h038A;
9'h19A: data = 16'h0001;
9'h19B: data = 16'h0000;
9'h19C: data = 16'h0380;
9'h19D: data = 16'h011C;
9'h19E: data = 16'h0000;
9'h19F: data = 16'h038A;
9'h1A0: data = 16'h0109;
9'h1A1: data = 16'h109C;
9'h1A2: data = 16'h0000;
9'h1A3: data = 16'h038A;
9'h1A4: data = 16'h0001;
9'h1A5: data = 16'h0000;
9'h1A6: data = 16'h0380;
9'h1A7: data = 16'h001C;
9'h1A8: data = 16'h0000;
9'h1A9: data = 16'h038E;
9'h1AA: data = 16'h002D;
9'h1AB: data = 16'h0000;
9'h1AC: data = 16'h00FF;
9'h1AD: data = 16'h0002;
9'h1AE: data = 16'h0000;
9'h1AF: data = 16'h01BC;
9'h1B0: data = 16'h001C;
9'h1B1: data = 16'h0000;
9'h1B2: data = 16'h038E;
9'h1B3: data = 16'h006D;
9'h1B4: data = 16'h0000;
9'h1B5: data = 16'h0008;
9'h1B6: data = 16'h0002;
9'h1B7: data = 16'h0000;
9'h1B8: data = 16'h01BC;
9'h1B9: data = 16'h011C;
9'h1BA: data = 16'h0000;
9'h1BB: data = 16'h038A;
9'h1BC: data = 16'h0109;
9'h1BD: data = 16'h109C;
9'h1BE: data = 16'h0000;
9'h1BF: data = 16'h038A;
9'h1C0: data = 16'h0370;
9'h1C1: data = 16'h0270;
9'h1C2: data = 16'h0170;
9'h1C3: data = 16'h0070;
9'h1C4: data = 16'h0090;
9'h1C5: data = 16'h0000;
9'h1C6: data = 16'h0000;
9'h1C7: data = 16'h0000;
9'h1C8: data = 16'h0000;
9'h1C9: data = 16'h0000;
9'h1CA: data = 16'h0000;
9'h1CB: data = 16'h0000;
9'h1CC: data = 16'hB000;
9'h1CD: data = 16'h0000;
9'h1CE: data = 16'h0000;
9'h1CF: data = 16'h0000;
9'h1D0: data = 16'h0000;
9'h1D1: data = 16'h0000;
9'h1D2: data = 16'h0000;


  endcase
endmodule
